library ieee;
use ieee.std_logic_1164.all;

entity  andN is
	generic (N : INTEGER  := 4); --bit  width
	port (
		A : in   std_logic_vector (N - 1  downto  0);
		B : in   std_logic_vector (N - 1  downto  0);
		Y : out  std_logic_vector (N - 1  downto  0)
	);
end  andN;

architecture generator of andN is
begin
	Y <= A and B;
end;
